sfkhdhsh
